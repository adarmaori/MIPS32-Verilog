module processor (
  input i_clk
);
  
endmodule
